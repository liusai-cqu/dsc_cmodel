package dsc_pkg;
  // 对应于C语言的枚举类型
  typedef enum int {
    FMT_RGB = 0,
    FMT_YUV = 1
  } format_t;
  
  typedef enum int {
    COLOR_RGB = 0,
    COLOR_YCC = 1
  } color_t;
  
  typedef enum int {
    CHROMA_444 = 0,
    CHROMA_422 = 1,
    CHROMA_420 = 2
  } chroma_t;
  
  typedef enum int {
    ALPHA_NONE = 0,
    ALPHA_USED = 1
  } alpha_t;
  
  // RGB数据结构
  typedef struct {
    int[][] r;
    int[][] g;
    int[][] b;
    int[][] a;
  } rgb_t;
  
  // YUV数据结构
  typedef struct {
    int[][] y;
    int[][] u;
    int[][] v;
  } yuv_t;
  
  // 图片数据联合体
  typedef union {
    rgb_t rgb;
    yuv_t yuv;
  } content_t;
  
  // 图片结构体
  typedef struct {
    format_t format;
    color_t color;
    chroma_t chroma;
    alpha_t alpha;
    int w;
    int h;
    int bits;
    int ar1;
    int ar2;
    int frm_no;
    int seq_len;
    real framerate;
    int interlaced;
    content_t data;
  } pic_t;
  
  // DSC配置结构体
  typedef struct {
    int slice_width;
    int slice_height;
    int bits_per_pixel;
    int bits_per_component;
    // 其他DSC配置参数
  } dsc_cfg_t;
  
  // 导入C函数的声明
  import "DPI-C" context function int dsc_algorithm_dpi(
    input int isEncoder,
    input dsc_cfg_t dsc_cfg,
    input pic_t ip,
    output pic_t op,
    inout byte unsigned cmpr_buf[],
    inout pic_t temp_pic[]
  );
  
endpackage : dsc_pkg
